** sch_path: /home/emman/Desktop/Acads/EE220/Simple-CS-Amplifier/csamp3.sch
**.subckt csamp3 vdd vdd vdd out
*.iopin vdd
*.iopin vdd
*.iopin vdd
*.opin out
XM1 net2 net1 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
E1 net1 GND net2 net3 1000
I0 vdd net2 3n
VDS net3 GND 0.9
V2 vdd GND 1.8
XM2 out in GND GND sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
I1 vdd out 3n
vin in net1 DC 0 AC 1
C1 out GND 5p m=1
**** begin user architecture code



.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.option wnflag=1 scale=1e-6

.control
save all

*save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[vgs]
*save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[vds]
*save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[gm]
*save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[id]
*save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[gds]
*save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cgg]

AC dec 10 1 100Meg

*let vgs = @m.xm2.msky130_fd_pr__nfet_01v8_lvt[vgs]
*let vds = @m.xm2.msky130_fd_pr__nfet_01v8_lvt[vds]
*let gm = @m.xm2.msky130_fd_pr__nfet_01v8_lvt[gm]
*let id = @m.xm2.msky130_fd_pr__nfet_01v8_lvt[id]
*let ro = 1/@m.xm2.msky130_fd_pr__nfet_01v8_lvt[gds]
*let cgg = @m.xm2.msky130_fd_pr__nfet_01v8_lvt[cgg]

*let ao = gm*ro
*let ft = gm/(2*pi*cgg)
*plot v(out)

*tran 10u 10m

*plot ao



*wrdata ao-L=0.40.txt ao
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
