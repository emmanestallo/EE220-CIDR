** sch_path: /home/emman/Desktop/Acads/EE220/Simple-CS-Amplifier/gmid.sch
**.subckt gmid
XM1 net2 net1 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
VGS net1 GND 0.9
VDS net2 GND 0.9
**** begin user architecture code



.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.option wnflag=1 scale=1e-6

.control

save all
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[id]
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gds]
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[w]
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cgg]
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vth]

dc VGS 0 1.8 1m

let id = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[id]
let gm = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
let ro = 1/@m.xm1.msky130_fd_pr__nfet_01v8_lvt[gds]
let width = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[w]
let cgg = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cgg]
let vth = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vth]

let gmoverid = gm/id
let vstar = 2/gmoverid
let gmro = gm*ro
let ft = gm/(2*pi*cgg)

*wrdata charac-L=0.23.txt ft gmro vstar

*meas dc gain find gmro when vstar=0.19
*meas dc freq find ft when vstar=0.19

*meas DC gain FIND gmro WHEN vstar=0.3
*meas DC freq FIND ft WHEN vstar=0.3
*meas DC current FIND id WHEN vstar=0.3

plot gmro



.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
