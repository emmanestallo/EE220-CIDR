** sch_path: /home/emman/Desktop/Acads/EE220/Simple-CS-Amplifier/csamp1.sch
**.subckt csamp1
XM1 net2 net1 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.40 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
E1 net1 GND net2 net4 1000
I0 net3 net2 1m
VDS net4 GND 1.8
V2 net3 GND 1.8
**** begin user architecture code



.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.option wnflag=1 scale=1e-6

.control
save all
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vgs]
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vds]
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gds]

dc VDS 0.2 1.8 1m

let vgs = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vgs]
let vds = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vds]
let gm = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
let gds = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gds]
let ro = 1/gds

let gain = gm*ro

let ao = -1/(deriv(vgs))

plot ao
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
