** sch_path: /home/emman/Desktop/Acads/EE220/MOS-Transition-Frequency/act5.sch
**.subckt act5 g1 d1
*.ipin g1
*.iopin d1
XM1 d1 g1 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.45 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.option wnflag = 1 scale=1e-6

vgs ga 0 dc=0.9
vds d1 0 dc=0.9

l1   ga g1 1e9
iac  g1 0 dc=0 ac=1
h1   io1 0 vds 1

.control
save all

save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[id]

let vgsx = 0
let run = 0
set curplot = new
set scratch = $curplot
let ft_vec = vector(181)
let vgs_vec = vector(181)

dowhile vgsx <= 1.81

  alter vgs = vgsx
  ac dec 100 1e6 1e12

  * plot vdb(io1)
  meas ac ft when vdb(io1) = 0

  set dt = $curplot
  setplot $scratch

  let vgs_vec[run] = vgsx
  let ft_vec[run] = {$dt}.ft

  setplot $dt

  echo Vgs {$&vgsx}
  echo ft {$&ft}
  echo Run {$&run}

  let vgsx = vgsx + 0.01
  let run = run + 1
end

setplot $scratch
setscale vgs_vec
wrdata mos-ft-tt-l=150nm-w=10um.dat ft_vec
plot ft_vec


.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
