** sch_path: /home/emman/Desktop/Acads/EE220/MOS-Design-Parameters/PMOS/act6.sch
**.subckt act6
XM1 net2 net1 GND GND sky130_fd_pr__pfet_01v8_lvt L=0.70 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
V1 GND net1 0.9
V2 GND net2 0.9
**** begin user architecture code



.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice ss
.option wnflag=1 scale=1e-6

.control

save all

save @m.xm1.msky130_fd_pr__pfet_01v8_lvt[id]
save @m.xm1.msky130_fd_pr__pfet_01v8_lvt[gm]


dc v1 -0.2 1.8 1m

let id = @m.xm1.msky130_fd_pr__pfet_01v8_lvt[id]
let gm = @m.xm1.msky130_fd_pr__pfet_01v8_lvt[gm]

let gmoverid = gm/id

#wrdata ftgmid-ss.txt ftgmid vstar

.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
