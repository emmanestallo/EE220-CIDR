** sch_path: /home/emman/Desktop/Acads/EE220/MOS-Transistor-Characteristics/act4p.sch
**.subckt act4p g1 d1
*.ipin g1
*.iopin d1
XM1 d1 g1 GND GND sky130_fd_pr__pfet_01v8_lvt L=1.05 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice ss
.option wnflag = 1 scale=1e-6

vgs g1 0 dc=-0.9
vds d1 0 dc=-0.9

.control
save all

save @m.xm1.msky130_fd_pr__pfet_01v8_lvt[id]

dc vgs 0 -1.8 -0.01
let idn = @m.xm1.msky130_fd_pr__pfet_01v8_lvt[id]
plot idn

wrdata mos-plvt-transfer-ss-l=1050nm-w=10um.dat idn

dc vds 0 -1.8 -0.01 vgs -0.45 -1.8 -0.45
let idn = @m.xm1.msky130_fd_pr__pfet_01v8_lvt[id]
plot idn

wrdata mos-plvt-output-ss-l=1050nm-w=10um.dat idn

.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
